library ieee;
use ieee.std_logic_1164.all;

-- Defining entities. Like a table of contents
entity example_and is
    port (
        input_1 : in std_logic;
        input_2 : in std_logic;
        and_result : out std_logic
        
    );
end example_and;


